/*a Copyright
  
  This file 'hierarchy_struct.cdl' copyright Gavin J Stark 2003, 2004
  
  This program is free software; you can redistribute it and/or modify it under
  the terms of the GNU General Public License as published by the Free Software
  Foundation, version 2.0.
  
  This program is distributed in the hope that it will be useful,
  but WITHOUT ANY WARRANTY; without even implied warranty of MERCHANTABILITY
  or FITNESS FOR A PARTICULAR PURPOSE. See the GNU General Public License
  for more details.
*/

/*a Includes
 */
include "test_hierarchy::hierarchy_struct.h"

/*a Module
 */
module hierarchy_struct( clock int_clock,
                         input bit int_reset,
                         input t_h_struct in,
                         output t_h_struct out )
{
    default clock int_clock;
    default reset int_reset;
    clocked t_h_struct out = { c=0, s={ x=0, y=0} };
    
    main_code "Main code":
        {
            out <= in;
        }
}

/*a Editor preferences and notes
mode: c ***
c-basic-offset: 4 ***
c-default-style: (quote ((c-mode . "k&r") (c++-mode . "k&r"))) ***
outline-regexp: "/\\\*a\\\|[\t ]*\/\\\*[b-z][\t ]" ***
*/

