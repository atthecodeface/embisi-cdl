/*a Copyright
  
  This file 'hierarchy_reg.cdl' copyright Gavin J Stark 2003, 2004
  
  This program is free software; you can redistribute it and/or modify it under
  the terms of the GNU General Public License as published by the Free Software
  Foundation, version 2.0.
  
  This program is distributed in the hope that it will be useful,
  but WITHOUT ANY WARRANTY; without even implied warranty of MERCHANTABILITY
  or FITNESS FOR A PARTICULAR PURPOSE. See the GNU General Public License
  for more details.
*/

/*a Includes
 */

/*a Module
 */
module hierarchy_reg2( clock int_clock,
                       clock int_bclock,
                       input bit int_reset,
                       input bit in,
                       output bit out,
    output bit out_b)
{
    default reset int_reset;
    clocked clock int_clock bit out = 0;
    clocked clock int_bclock bit out_b = 0;

    main_code "Main code":
        {
            out <= in;
            out_b <= in;
        }
}

/*a Editor preferences and notes
mode: c ***
c-basic-offset: 4 ***
c-default-style: (quote ((c-mode . "k&r") (c++-mode . "k&r"))) ***
outline-regexp: "/\\\*a\\\|[\t ]*\/\\\*[b-z][\t ]" ***
*/

